***********************************************************
*
* BCV26
*
* Nexperia
*
* Darlington PNP Transistor
* IC   = 500 mA
* VCEO = 30 V 
* hFE  = min 20000 @ 5V/100mA
* 
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base  
* Package Pin 2: Emitter
* Package Pin 3: Collector
* 
*
* # 
* Spicemodel does not include temperature dependency
*
**********************************************************
*#
*
* For use with Microsim PSPICE 
* please modify the AREA statement
* in this model:  e.g.
* SPICE: 
* Q2 3 22 2 BCV26 AREA = 4.68 
* PSPICE:
* Q2 3 22 2 BCV26 4.68 
*
.SUBCKT BCV26 1 2 3
Q1 1 2 33 BCV26 1 
Q2 1 33 3 BCV26 4.68
*
.MODEL BCV26 PNP 
+ IS = 1.593E-14 
+ NF = 0.9855 
+ ISE = 7E-15 
+ NE = 1.5 
+ BF = 280 
+ IKF = 0.09 
+ VAF = 31 
+ NR = 1 
+ ISC = 1E-32 
+ NC = 2 
+ BR = 5 
+ IKR = 0.1 
+ VAR = 4 
+ RB = 600 
+ IRB = 1E-06 
+ RBM = 10 
+ RE = 0.1 
+ RC = 1 
+ XTB = 0 
+ EG = 1.11 
+ XTI = 3 
+ CJE = 1.32E-11 
+ VJE = 0.9 
+ MJE = 0.4141 
+ TF = 9.9E-10 
+ XTF = 15 
+ VTF = 5 
+ ITF = 0.4 
+ PTF = 0 
+ CJC = 7.95E-12 
+ VJC = 0.9 
+ MJC = 0.5622 
+ XCJC = 0.9 
+ TR = 1E-15 
+ CJS = 0 
+ VJS = 0.75 
+ MJS = 0.333 
+ FC = 0.98
.ENDS
*