***********************************************************
*
* BCV27
*
* Nexperia
*
* Darlington NPN Transistor
* IC   = 500 mA
* VCEO = 30 V 
* hFE  = 20000 @ 5V/100mA
* 
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base  
* Package Pin 2: Emitter
* Package Pin 3: Collector
* 
*
* # 
* Spicemodel does not include temperature dependency
*
**********************************************************
*#
*
* For use with Microsim PSPICE 
* please modify the AREA statement
* in this model:  e.g.
* SPICE: 
* Q2 3 22 2 BCV27 AREA = 5.1 
* PSPICE:
* Q2 3 22 2 BCV27 5.1 
* VTF, ITF, XTF are set to 
* default values 
*
.SUBCKT BCV27 1 2 3
Q1 1 2 33 BCV27 1 
Q2 1 33 3 BCV27 5.1 
*
.MODEL BCV27 NPN 
+ IS = 1.35E-14 
+ NF = 0.9889 
+ ISE = 4.441E-28 
+ NE = 1.03 
+ BF = 204 
+ IKF = 0.1 
+ VAF = 94 
+ NR = 1 
+ ISC = 1E-32 
+ NC = 2 
+ BR = 5 
+ IKR = 0.1 
+ VAR = 10 
+ RB = 45 
+ IRB = 7E-06 
+ RBM = 1 
+ RE = 0.25 
+ RC = 2 
+ XTB = 0 
+ EG = 1.11 
+ XTI = 3 
+ CJE = 1.445E-11 
+ VJE = 0.9 
+ MJE = 0.3635 
+ TF = 7E-10 
+ XTF = 1 
+ VTF = 1000 
+ ITF = 0.01 
+ PTF = 0 
+ CJC = 4.89E-12 
+ VJC = 0.6559 
+ MJC = 0.5115 
+ XCJC = 1 
+ TR = 1E-07 
+ CJS = 0 
+ VJS = 0.75 
+ MJS = 0.333 
+ FC = 0.999 
.ENDS
*